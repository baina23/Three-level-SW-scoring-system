`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/08/20 10:45:29
// Design Name: 
// Module Name: SW
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SW(
input clk,
input rst,
input [71:0] ref,
input [71:0] read,
output reg[6:0] max,
output [12:0] loc,
output reg finish
    );
parameter l = 16;
reg [6:0] state;
reg[12:0] loc1,loc2;
reg[1:0] sig;
reg rst1;

wire [6:0] d1_01, d1_02, d1_10,d1_20,d1_3;
wire [6:0] d2_01, d2_02, d2_10,d2_20,d2_3;
wire [6:0] d3_01, d3_02, d3_10,d3_20,d3_3;
wire [6:0] d4_01, d4_02, d4_10,d4_20,d4_3;
wire [6:0] d5_01, d5_02, d5_10,d5_20,d5_3;
wire [6:0] d6_01, d6_02, d6_10,d6_20,d6_3;
wire [6:0] d7_01, d7_02, d7_10,d7_20,d7_3;
wire [6:0] d8_01, d8_02, d8_10,d8_20,d8_3;
wire [6:0] d9_01, d9_02, d9_10,d9_20,d9_3;
wire [6:0] d10_01, d10_02, d10_10,d10_20,d10_3;
wire [6:0] d11_01, d11_02, d11_10,d11_20,d11_3;
wire [6:0] d12_01, d12_02, d12_10,d12_20,d12_3;

reg [6:0] D1_3, DD1_3, DDD1_3;//, DDDD1_3, DDDDD1_3, DDDDDD1_3;
reg [6:0] D2_3, DD2_3, DDD2_3;//, DDDD2_3, DDDDD2_3, DDDDDD2_3;
reg [6:0] D3_3, DD3_3, DDD3_3;//, DDDD3_3, DDDDD3_3, DDDDDD3_3;
reg [6:0] D4_3, DD4_3, DDD4_3;//, DDDD4_3, DDDDD4_3, DDDDDD4_3;
reg [6:0] D5_3, DD5_3, DDD5_3;//, DDDD5_3, DDDDD5_3, DDDDDD5_3;
reg [6:0] D6_3, DD6_3, DDD6_3;//, DDDD6_3, DDDDD6_3, DDDDDD6_3;
reg [6:0] D7_3, DD7_3, DDD7_3;//, DDDD7_3, DDDDD7_3, DDDDDD7_3;
reg [6:0] D8_3, DD8_3, DDD8_3;//, DDDD8_3, DDDDD8_3, DDDDDD8_3;
reg [6:0] D9_3, DD9_3, DDD9_3;//, DDDD9_3, DDDDD9_3, DDDDDD9_3;
reg [6:0] D10_3, DD10_3, DDD10_3;//, DDDD10_3, DDDDD10_3, DDDDDD10_3;
reg [6:0] D11_3, DD11_3, DDD11_3;//, DDDD11_3, DDDDD11_3, DDDDDD11_3;
reg [6:0] D12_3, DD12_3, DDD12_3;//, DDDD12_3, DDDDD12_3, DDDDDD12_3;


reg [5:0] seq_1,targ_1;
reg[6:0] f00_1,f01_1,f02_1,f03_1,f10_1,f20_1,f30_1;
wire[6:0] f11_1,f12_1,f13_1,f21_1,f22_1,f23_1,f31_1,f32_1,f33_1;
//wire[6:0] F11_1,F12_1,F13_1,F21_1,F22_1,F23_1,F31_1,F32_1,F33_1;

reg [5:0] seq_2,targ_2;
reg[6:0] f00_2,f01_2,f02_2,f03_2,f10_2,f20_2,f30_2;
wire[6:0] f11_2,f12_2,f13_2,f21_2,f22_2,f23_2,f31_2,f32_2,f33_2;
//wire[6:0] F11_2,F12_2,F13_2,F21_2,F22_2,F23_2,F31_2,F32_2,F33_2;

reg [5:0] seq_3,targ_3;
reg[6:0] f00_3,f01_3,f02_3,f03_3,f10_3,f20_3,f30_3;
wire[6:0] f11_3,f12_3,f13_3,f21_3,f22_3,f23_3,f31_3,f32_3,f33_3;
//wire[6:0] F11_3,F12_3,F13_3,F21_3,F22_3,F23_3,F31_3,F32_3,F33_3;

reg [5:0] seq_4,targ_4;
reg[6:0] f00_4,f01_4,f02_4,f03_4,f10_4,f20_4,f30_4;
wire[6:0] f11_4,f12_4,f13_4,f21_4,f22_4,f23_4,f31_4,f32_4,f33_4;
//wire[6:0] F11_4,F12_4,F13_4,F21_4,F22_4,F23_4,F31_4,F32_4,F33_4;

reg [5:0] seq_5,targ_5;
reg[6:0] f00_5,f01_5,f02_5,f03_5,f10_5,f20_5,f30_5;
wire[6:0] f11_5,f12_5,f13_5,f21_5,f22_5,f23_5,f31_5,f32_5,f33_5;
//wire[6:0] F11_5,F12_5,F13_5,F21_5,F22_5,F23_5,F31_5,F32_5,F33_5;

reg [5:0] seq_6,targ_6;
reg[6:0] f00_6,f01_6,f02_6,f03_6,f10_6,f20_6,f30_6;
wire[6:0] f11_6,f12_6,f13_6,f21_6,f22_6,f23_6,f31_6,f32_6,f33_6;
//wire[6:0]F11_6,F12_6,F13_6,F21_6,F22_6,F23_6,F31_6,F32_6,F33_6;

reg [5:0] seq_7,targ_7;
reg[6:0] f00_7,f01_7,f02_7,f03_7,f10_7,f20_7,f30_7;
wire[6:0] f11_7,f12_7,f13_7,f21_7,f22_7,f23_7,f31_7,f32_7,f33_7;
//wire[6:0]F11_7,F12_7,F13_7,F21_7,F22_7,F23_7,F31_7,F32_7,F33_7;

reg [5:0] seq_8,targ_8;
reg[6:0] f00_8,f01_8,f02_8,f03_8,f10_8,f20_8,f30_8;
wire[6:0] f11_8,f12_8,f13_8,f21_8,f22_8,f23_8,f31_8,f32_8,f33_8;
//wire[6:0]F11_8,F12_8,F13_8,F21_8,F22_8,F23_8,F31_8,F32_8,F33_8;

reg [5:0] seq_9,targ_9;
reg[6:0] f00_9,f01_9,f02_9,f03_9,f10_9,f20_9,f30_9;
wire[6:0] f11_9,f12_9,f13_9,f21_9,f22_9,f23_9,f31_9,f32_9,f33_9;
//wire[6:0]F11_9,F12_9,F13_9,F21_9,F22_9,F23_9,F31_9,F32_9,F33_9;

reg [5:0] seq_10,targ_10;
reg[6:0] f00_10,f01_10,f02_10,f03_10,f10_10,f20_10,f30_10;
wire[6:0] f11_10,f12_10,f13_10,f21_10,f22_10,f23_10,f31_10,f32_10,f33_10;
//wire[6:0]F11_10,F12_10,F13_10,F21_10,F22_10,F23_10,F31_10,F32_10,F33_10;

reg [5:0] seq_11,targ_11;
reg[6:0] f00_11,f01_11,f02_11,f03_11,f10_11,f20_11,f30_11;
wire[6:0] f11_11,f12_11,f13_11,f21_11,f22_11,f23_11,f31_11,f32_11,f33_11;
//wire[6:0]F11_11,F12_11,F13_11,F21_11,F22_11,F23_11,F31_11,F32_11,F33_11;

reg [5:0] seq_12,targ_12;
reg[6:0] f00_12,f01_12,f02_12,f03_12,f10_12,f20_12,f30_12;
wire[6:0] f11_12,f12_12,f13_12,f21_12,f22_12,f23_12,f31_12,f32_12,f33_12;
//wire[6:0]F11_12,F12_12,F13_12,F21_12,F22_12,F23_12,F31_12,F32_12,F33_12;



SW_core PE1(.clk(clk),.rst(rst1),.seq(seq_1),.targ(targ_1),.f00(f00_1),.f01(f01_1),.f02(f02_1),.f03(f03_1),.f10(f10_1),.f20(f20_1),.f30(f30_1),.f11(f11_1),.f12(f12_1),.f13(f13_1),.f21(f21_1),.f22(f22_1),.f23(f23_1),.f31(f31_1),.f32(f32_1),.f33(f33_1) );
SW_core PE2(.clk(clk),.rst(rst1),.seq(seq_2),.targ(targ_2),.f00(f00_2),.f01(f01_2),.f02(f02_2),.f03(f03_2),.f10(f10_2),.f20(f20_2),.f30(f30_2),.f11(f11_2),.f12(f12_2),.f13(f13_2),.f21(f21_2),.f22(f22_2),.f23(f23_2),.f31(f31_2),.f32(f32_2),.f33(f33_2));
SW_core PE3(.clk(clk),.rst(rst1),.seq(seq_3),.targ(targ_3),.f00(f00_3),.f01(f01_3),.f02(f02_3),.f03(f03_3),.f10(f10_3),.f20(f20_3),.f30(f30_3),.f11(f11_3),.f12(f12_3),.f13(f13_3),.f21(f21_3),.f22(f22_3),.f23(f23_3),.f31(f31_3),.f32(f32_3),.f33(f33_3) );
SW_core PE4(.clk(clk),.rst(rst1),.seq(seq_4),.targ(targ_4),.f00(f00_4),.f01(f01_4),.f02(f02_4),.f03(f03_4),.f10(f10_4),.f20(f20_4),.f30(f30_4),.f11(f11_4),.f12(f12_4),.f13(f13_4),.f21(f21_4),.f22(f22_4),.f23(f23_4),.f31(f31_4),.f32(f32_4),.f33(f33_4) );
SW_core PE5(.clk(clk),.rst(rst1),.seq(seq_5),.targ(targ_5),.f00(f00_5),.f01(f01_5),.f02(f02_5),.f03(f03_5),.f10(f10_5),.f20(f20_5),.f30(f30_5),.f11(f11_5),.f12(f12_5),.f13(f13_5),.f21(f21_5),.f22(f22_5),.f23(f23_5),.f31(f31_5),.f32(f32_5),.f33(f33_5) );
SW_core PE6(.clk(clk),.rst(rst1),.seq(seq_6),.targ(targ_6),.f00(f00_6),.f01(f01_6),.f02(f02_6),.f03(f03_6),.f10(f10_6),.f20(f20_6),.f30(f30_6),.f11(f11_6),.f12(f12_6),.f13(f13_6),.f21(f21_6),.f22(f22_6),.f23(f23_6),.f31(f31_6),.f32(f32_6),.f33(f33_6) );
SW_core PE7(.clk(clk),.rst(rst1),.seq(seq_7),.targ(targ_7),.f00(f00_7),.f01(f01_7),.f02(f02_7),.f03(f03_7),.f10(f10_7),.f20(f20_7),.f30(f30_7),.f11(f11_7),.f12(f12_7),.f13(f13_7),.f21(f21_7),.f22(f22_7),.f23(f23_7),.f31(f31_7),.f32(f32_7),.f33(f33_7) );
SW_core PE8(.clk(clk),.rst(rst1),.seq(seq_8),.targ(targ_8),.f00(f00_8),.f01(f01_8),.f02(f02_8),.f03(f03_8),.f10(f10_8),.f20(f20_8),.f30(f30_8),.f11(f11_8),.f12(f12_8),.f13(f13_8),.f21(f21_8),.f22(f22_8),.f23(f23_8),.f31(f31_8),.f32(f32_8),.f33(f33_8) );
SW_core PE9(.clk(clk),.rst(rst1),.seq(seq_9),.targ(targ_9),.f00(f00_9),.f01(f01_9),.f02(f02_9),.f03(f03_9),.f10(f10_9),.f20(f20_9),.f30(f30_9),.f11(f11_9),.f12(f12_9),.f13(f13_9),.f21(f21_9),.f22(f22_9),.f23(f23_9),.f31(f31_9),.f32(f32_9),.f33(f33_9) );
SW_core PE10(.clk(clk),.rst(rst1),.seq(seq_10),.targ(targ_10),.f00(f00_10),.f01(f01_10),.f02(f02_10),.f03(f03_10),.f10(f10_10),.f20(f20_10),.f30(f30_10),.f11(f11_10),.f12(f12_10),.f13(f13_10),.f21(f21_10),.f22(f22_10),.f23(f23_10),.f31(f31_10),.f32(f32_10),.f33(f33_10) );
SW_core PE11(.clk(clk),.rst(rst1),.seq(seq_11),.targ(targ_11),.f00(f00_11),.f01(f01_11),.f02(f02_11),.f03(f03_11),.f10(f10_11),.f20(f20_11),.f30(f30_11),.f11(f11_11),.f12(f12_11),.f13(f13_11),.f21(f21_11),.f22(f22_11),.f23(f23_11),.f31(f31_11),.f32(f32_11),.f33(f33_11) );
SW_core PE12(.clk(clk),.rst(rst1),.seq(seq_12),.targ(targ_12),.f00(f00_12),.f01(f01_12),.f02(f02_12),.f03(f03_12),.f10(f10_12),.f20(f20_12),.f30(f30_12),.f11(f11_12),.f12(f12_12),.f13(f13_12),.f21(f21_12),.f22(f22_12),.f23(f23_12),.f31(f31_12),.f32(f32_12),.f33(f33_12) );


assign d1_01 = f31_1; 
assign d1_02 = f32_1;
assign d1_10 = f13_1;
assign d1_20 = f23_1;
assign d1_3 = f33_1;
assign d2_01 = f31_2;
assign d2_02 = f32_2;
assign d2_10 = f13_2;
assign d2_20 = f23_2;
assign d2_3 = f33_2; 
assign d3_01 = f31_3;
assign d3_02 = f32_3;
assign d3_10 = f13_3;
assign d3_20 = f23_3;
assign d3_3 = f33_3;
assign d4_01 = f31_4;
assign d4_02 = f32_4;
assign d4_10 = f13_4;
assign d4_20 = f23_4;
assign d4_3 = f33_4;
assign d5_01 = f31_5;
assign d5_02 = f32_5;
assign d5_10 = f13_5;
assign d5_20 = f23_5;
assign d5_3 = f33_5;
assign d6_01 = f31_6;
assign d6_02 = f32_6;
assign d6_10 = f13_6;
assign d6_20 = f23_6;
assign d6_3 = f33_6;
assign d7_01 = f31_7;
assign d7_02 = f32_7;
assign d7_10 = f13_7;
assign d7_20 = f23_7;
assign d7_3 = f33_7;
assign d8_01 = f31_8;
assign d8_02 = f32_8;
assign d8_10 = f13_8;
assign d8_20 = f23_8;
assign d8_3 = f33_8;
assign d9_01 = f31_9;
assign d9_02 = f32_9;
assign d9_10 = f13_9;
assign d9_20 = f23_9;
assign d9_3 = f33_9;
assign d10_01 = f31_10;
assign d10_02 = f32_10;
assign d10_10 = f13_10;
assign d10_20 = f23_10;
assign d10_3 = f33_10;
assign d11_01 = f31_11;
assign d11_02 = f32_11;
assign d11_10 = f13_11;
assign d11_20 = f23_11;
assign d11_3 = f33_11;
assign d12_01 = f31_12;
assign d12_02 = f32_12;
assign d12_10 = f13_12;
assign d12_20 = f23_12;
assign d12_3 = f33_12;

assign loc = (sig == 2'b00)?13'd0:
             (sig == 2'b01)?loc1:
             (sig == 2'b10)?loc2:
             (sig == 2'b11)?(loc1|loc2):13'd0;


always@(posedge clk)
begin
    if(!rst)
        begin
        state <= 0;
        rst1 <= 0;
        max <= 5'd0;
        loc1 <= 13'd0;
        loc2 <= 13'd0;
        sig <= 2'b00;
        finish <= 1;
        seq_1 <= 6'b000000;targ_1 <= 6'b111111;f00_1 <= l;f01_1 <= l;f02_1 <= l;f03_1 <= l;f10_1 <= l;f20_1 <= l;f30_1 <= l;
        seq_2 <= 6'b000000;targ_2 <= 6'b111111;f00_2 <= l;f01_2 <= l;f02_2 <= l;f03_2 <= l;f10_2 <= l;f20_2 <= l;f30_2 <= l;
        seq_3 <= 6'b000000;targ_3 <= 6'b111111;f00_3 <= l;f01_3 <= l;f02_3 <= l;f03_3 <= l;f10_3 <= l;f20_3 <= l;f30_3 <= l;
        seq_4 <= 6'b000000;targ_4 <= 6'b111111;f00_4 <= l;f01_4 <= l;f02_4 <= l;f03_4 <= l;f10_4 <= l;f20_4 <= l;f30_4 <= l;
        seq_5 <= 6'b000000;targ_5 <= 6'b111111;f00_5 <= l;f01_5 <= l;f02_5 <= l;f03_5 <= l;f10_5 <= l;f20_5 <= l;f30_5 <= l;
        seq_6 <= 6'b000000;targ_6 <= 6'b111111;f00_6 <= l;f01_6 <= l;f02_6 <= l;f03_6 <= l;f10_6 <= l;f20_6 <= l;f30_6 <= l;
        seq_7 <= 6'b000000;targ_7 <= 6'b111111;f00_7 <= l;f01_7 <= l;f02_7 <= l;f03_7 <= l;f10_7 <= l;f20_7 <= l;f30_7 <= l;
        seq_8 <= 6'b000000;targ_8 <= 6'b111111;f00_8 <= l;f01_8 <= l;f02_8 <= l;f03_8 <= l;f10_8 <= l;f20_8 <= l;f30_8 <= l;
        seq_9 <= 6'b000000;targ_9 <= 6'b111111;f00_9 <= l;f01_9 <= l;f02_9 <= l;f03_9 <= l;f10_9 <= l;f20_9 <= l;f30_9 <= l;
        seq_10 <= 6'b000000;targ_10 <= 6'b111111;f00_10 <= l;f01_10 <= l;f02_10 <= l;f03_10 <= l;f10_10 <= l;f20_10 <= l;f30_10 <= l;
        seq_11 <= 6'b000000;targ_11 <= 6'b111111;f00_11 <= l;f01_11 <= l;f02_11 <= l;f03_11 <= l;f10_11 <= l;f20_11 <= l;f30_11 <= l;      
        seq_12 <= 6'b000000;targ_12 <= 6'b111111;f00_12 <= l;f01_12 <= l;f02_12 <= l;f03_12 <= l;f10_12 <= l;f20_12 <= l;f30_12 <= l;            
       
        D1_3 <= 0;
        D2_3 <= 0;
        D3_3 <= 0;
        D4_3 <= 0;
        D5_3 <= 0;
        D6_3 <= 0;
        D7_3 <= 0;
        D8_3 <= 0;
        D9_3 <= 0;
        D10_3 <= 0;
        D11_3 <= 0;
        D12_3 <= 0;  
       
       end
   
    else 
    begin
        D1_3 <= DD1_3;DD1_3 <=  DDD1_3;DDD1_3 <= d1_3;//DDDD1_3;DDDD1_3 <= DDDDD1_3;DDDDD1_3 <= DDDDDD1_3;DDDDDD1_3 <= d1_3;
        D2_3 <= DD2_3;DD2_3 <=  DDD2_3;DDD2_3 <= d2_3;//DDDD2_3;DDDD2_3 <= DDDDD2_3;DDDDD2_3 <= DDDDDD1_3;DDDDDD2_3 <= d2_3;
        D3_3 <= DD3_3;DD3_3 <= DDD3_3;DDD3_3 <= d3_3;//DDDD3_3;DDDD3_3 <= DDDDD3_3;DDDDD3_3 <= DDDDDD1_3;DDDDDD3_3 <= d3_3;
        D4_3 <= DD4_3;DD4_3 <= DDD4_3;DDD4_3 <= d4_3;//DDDD4_3;DDDD4_3 <= DDDDD4_3;DDDDD4_3 <= DDDDDD1_3;DDDDDD4_3 <= d4_3;
        D5_3 <= DD5_3;DD5_3 <= DDD5_3;DDD5_3 <= d5_3;//DDDD5_3;DDDD5_3 <= DDDDD5_3;DDDDD5_3 <= DDDDDD1_3;DDDDDD5_3 <= d5_3;
        D6_3 <= DD6_3;DD6_3 <= DDD6_3;DDD6_3 <= d6_3;//DDDD6_3;DDDD6_3 <= DDDDD6_3;DDDDD6_3 <= DDDDDD1_3;DDDDDD6_3 <= d6_3;
        D7_3 <= DD7_3;DD7_3 <= DDD7_3;DDD7_3 <= d7_3;//DDDD7_3;DDDD7_3 <= DDDDD7_3;DDDDD7_3 <= DDDDDD1_3;DDDDDD7_3 <= d7_3;
        D8_3 <= DD8_3;DD8_3 <= DDD8_3;DDD8_3 <= d8_3;//DDDD8_3;DDDD8_3 <= DDDDD8_3;DDDDD8_3 <= DDDDDD1_3;DDDDDD8_3 <= d8_3;
        D9_3 <= DD9_3;DD9_3 <= DDD9_3;DDD9_3 <= d9_3;//DDDD9_3;DDDD9_3 <= DDDDD9_3;DDDDD9_3 <= DDDDDD1_3;DDDDDD9_3 <= d9_3;
        D10_3 <= DD10_3;DD10_3 <= DDD10_3;DDD10_3 <= d10_3;//DDDD10_3;DDDD10_3 <= DDDDD10_3;DDDDD10_3 <= DDDDDD1_3;DDDDDD10_3 <= d10_3;
        D11_3 <= DD11_3;DD11_3 <= DDD11_3;DDD11_3 <= d11_3;//DDDD11_3;DDDD11_3 <= DDDDD11_3;DDDDD11_3 <= DDDDDD1_3;DDDDDD11_3 <= d11_3;
        D12_3 <= DD12_3;DD12_3 <= DDD12_3;DDD12_3 <= d12_3;//DDDD12_3;DDDD12_3 <= DDDDD12_3;DDDDD12_3 <= DDDDDD1_3;DDDDDD12_3 <= d12_3;
        finish <= 0;      
    case(state)
        7'd0:begin
                state <= state + 1;
                rst1 <= 1;
             end
        7'd1:
            begin
                seq_1 <= ref[71:66];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= l;f02_1 <= l;f03_1 <= l;f10_1 <= l;f20_1 <= l;f30_1 <= l;          
                state <= state + 1;                
            end
        7'd4:
            begin
                seq_1 <= ref[65:60];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= d1_01;f02_1 <= d1_02;f03_1 <= d1_3;f10_1 <= l;f20_1 <= l;f30_1 <= l;
                seq_2 <= ref[71:66];targ_2 <= read[65:60];f00_2 <= l;f01_2 <= l;f02_2 <= l;f03_2 <= l;f10_2 <= d1_10;f20_2 <= d1_20;f30_2 <= d1_3;               
                state <= state + 1;
            end 
        7'd7:
            begin
                seq_1 <= ref[59:54];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= d1_01;f02_1 <= d1_02;f03_1 <= d1_3;f10_1 <= l;f20_1 <= l;f30_1 <= l;
                seq_2 <= ref[65:60];targ_2 <= read[65:60];f00_2 <= D1_3;f01_2 <= d2_01;f02_2 <= d2_02;f03_2 <= d2_3;f10_2 <= d1_10;f20_2 <= d1_20;f30_2 <= d1_3;     
                seq_3 <= ref[71:66];targ_3 <= read[59:54];f00_3 <= l;f01_3 <= l;f02_3 <= l;f03_3 <= l;f10_3 <= d2_10;f20_3 <= d2_20;f30_3 <= d2_3;
                state <= state + 1;
             end
        7'd10:
            begin
                seq_1 <= ref[53:48];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= d1_01;f02_1 <= d1_02;f03_1 <= d1_3;f10_1 <= l;f20_1 <= l;f30_1 <= l;
                seq_2 <= ref[59:54];targ_2 <= read[65:60];f00_2 <= D1_3;f01_2 <= d2_01;f02_2 <= d2_02;f03_2 <= d2_3;f10_2 <= d1_10;f20_2 <= d1_20;f30_2 <= d1_3;
                seq_3 <= ref[65:60];targ_3 <= read[59:54];f00_3 <= D2_3;f01_3 <= d3_01;f02_3 <= d3_02;f03_3 <= d3_3;f10_3 <= d2_10;f20_3 <= d2_20;f30_3 <= d2_3;     
                seq_4 <= ref[71:66];targ_4 <= read[53:48];f00_4 <= l;f01_4 <= l;f02_4 <= l;f03_4 <= l;f10_4 <= d3_10;f20_4 <= d3_20;f30_4 <= d3_3;
                state <= state + 1;
            end
       7'd13:
            begin
                seq_1 <= ref[47:42];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= d1_01;f02_1 <= d1_02;f03_1 <= d1_3;f10_1 <= l;f20_1 <= l;f30_1 <= l;
                seq_2 <= ref[53:48];targ_2 <= read[65:60];f00_2 <= D1_3;f01_2 <= d2_01;f02_2 <= d2_02;f03_2 <= d2_3;f10_2 <= d1_10;f20_2 <= d1_20;f30_2 <= d1_3;
                seq_3 <= ref[59:54];targ_3 <= read[59:54];f00_3 <= D2_3;f01_3 <= d3_01;f02_3 <= d3_02;f03_3 <= d3_3;f10_3 <= d2_10;f20_3 <= d2_20;f30_3 <= d2_3;
                seq_4 <= ref[65:60];targ_4 <= read[53:48];f00_4 <= D3_3;f01_4 <= d4_01;f02_4 <= d4_02;f03_4 <= d4_3;f10_4 <= d3_10;f20_4 <= d3_20;f30_4 <= d3_3;     
                seq_5 <= ref[71:66];targ_5 <= read[47:42];f00_5 <= l;f01_5 <= l;f02_5 <= l;f03_5 <= l;f10_5 <= d4_10;f20_5 <= d4_20;f30_5 <= d4_3;
                state <= state + 1;
            end
       7'd16:
            begin
                seq_1 <= ref[41:36];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= d1_01;f02_1 <= d1_02;f03_1 <= d1_3;f10_1 <= l;f20_1 <= l;f30_1 <= l;
                seq_2 <= ref[47:42];targ_2 <= read[65:60];f00_2 <= D1_3;f01_2 <= d2_01;f02_2 <= d2_02;f03_2 <= d2_3;f10_2 <= d1_10;f20_2 <= d1_20;f30_2 <= d1_3;
                seq_3 <= ref[53:48];targ_3 <= read[59:54];f00_3 <= D2_3;f01_3 <= d3_01;f02_3 <= d3_02;f03_3 <= d3_3;f10_3 <= d2_10;f20_3 <= d2_20;f30_3 <= d2_3;
                seq_4 <= ref[59:54];targ_4 <= read[53:48];f00_4 <= D3_3;f01_4 <= d4_01;f02_4 <= d4_02;f03_4 <= d4_3;f10_4 <= d3_10;f20_4 <= d3_20;f30_4 <= d3_3;     
                seq_5 <= ref[65:60];targ_5 <= read[47:42];f00_5 <= D4_3;f01_5 <= d5_01;f02_5 <= d5_02;f03_5 <= d5_3;f10_5 <= d4_10;f20_5 <= d4_20;f30_5 <= d4_3;
                seq_6 <= ref[71:66];targ_6 <= read[41:36];f00_6 <= l;f01_6 <= l;f02_6 <= l;f03_6 <= l;f10_6 <= d5_10;f20_6 <= d5_20;f30_6 <= d5_3;
                state <= state + 1;
            end
       7'd19:
            begin
                seq_1 <= ref[35:30];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= d1_01;f02_1 <= d1_02;f03_1 <= d1_3;f10_1 <= l;f20_1 <= l;f30_1 <= l;
                seq_2 <= ref[41:36];targ_2 <= read[65:60];f00_2 <= D1_3;f01_2 <= d2_01;f02_2 <= d2_02;f03_2 <= d2_3;f10_2 <= d1_10;f20_2 <= d1_20;f30_2 <= d1_3;
                seq_3 <= ref[47:42];targ_3 <= read[59:54];f00_3 <= D2_3;f01_3 <= d3_01;f02_3 <= d3_02;f03_3 <= d3_3;f10_3 <= d2_10;f20_3 <= d2_20;f30_3 <= d2_3;
                seq_4 <= ref[53:48];targ_4 <= read[53:48];f00_4 <= D3_3;f01_4 <= d4_01;f02_4 <= d4_02;f03_4 <= d4_3;f10_4 <= d3_10;f20_4 <= d3_20;f30_4 <= d3_3;     
                seq_5 <= ref[59:54];targ_5 <= read[47:42];f00_5 <= D4_3;f01_5 <= d5_01;f02_5 <= d5_02;f03_5 <= d5_3;f10_5 <= d4_10;f20_5 <= d4_20;f30_5 <= d4_3;
                seq_6 <= ref[65:60];targ_6 <= read[41:36];f00_6 <= D5_3;f01_6 <= d6_01;f02_6 <= d6_02;f03_6 <= d6_3;f10_6 <= d5_10;f20_6 <= d5_20;f30_6 <= d5_3;
                seq_7 <= ref[71:66];targ_7 <= read[35:30];f00_7 <= l;f01_7 <= l;f02_7 <= l;f03_7 <= l;f10_7 <= d6_10;f20_7 <= d6_20;f30_7 <= d6_3;
                state <= state + 1;
            end
       7'd22:
            begin
                seq_1 <= ref[29:24];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= d1_01;f02_1 <= d1_02;f03_1 <= d1_3;f10_1 <= l;f20_1 <= l;f30_1 <= l;
                seq_2 <= ref[35:30];targ_2 <= read[65:60];f00_2 <= D1_3;f01_2 <= d2_01;f02_2 <= d2_02;f03_2 <= d2_3;f10_2 <= d1_10;f20_2 <= d1_20;f30_2 <= d1_3;
                seq_3 <= ref[41:36];targ_3 <= read[59:54];f00_3 <= D2_3;f01_3 <= d3_01;f02_3 <= d3_02;f03_3 <= d3_3;f10_3 <= d2_10;f20_3 <= d2_20;f30_3 <= d2_3;
                seq_4 <= ref[47:42];targ_4 <= read[53:48];f00_4 <= D3_3;f01_4 <= d4_01;f02_4 <= d4_02;f03_4 <= d4_3;f10_4 <= d3_10;f20_4 <= d3_20;f30_4 <= d3_3;     
                seq_5 <= ref[53:48];targ_5 <= read[47:42];f00_5 <= D4_3;f01_5 <= d5_01;f02_5 <= d5_02;f03_5 <= d5_3;f10_5 <= d4_10;f20_5 <= d4_20;f30_5 <= d4_3;
                seq_6 <= ref[59:54];targ_6 <= read[41:36];f00_6 <= D5_3;f01_6 <= d6_01;f02_6 <= d6_02;f03_6 <= d6_3;f10_6 <= d5_10;f20_6 <= d5_20;f30_6 <= d5_3;
                seq_7 <= ref[65:60];targ_7 <= read[35:30];f00_7 <= D6_3;f01_7 <= d7_01;f02_7 <= d7_02;f03_7 <= d7_3;f10_7 <= d6_10;f20_7 <= d6_20;f30_7 <= d6_3;
                seq_8 <= ref[71:66];targ_8 <= read[29:24];f00_8 <= l;f01_8 <= l;f02_8 <= l;f03_8 <= l;f10_8 <= d7_10;f20_8 <= d7_20;f30_8 <= d7_3;
                state <= state + 1;
            end
       7'd25:
            begin
                seq_1 <= ref[23:18];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= d1_01;f02_1 <= d1_02;f03_1 <= d1_3;f10_1 <= l;f20_1 <= l;f30_1 <= l;
                seq_2 <= ref[29:24];targ_2 <= read[65:60];f00_2 <= D1_3;f01_2 <= d2_01;f02_2 <= d2_02;f03_2 <= d2_3;f10_2 <= d1_10;f20_2 <= d1_20;f30_2 <= d1_3;
                seq_3 <= ref[35:30];targ_3 <= read[59:54];f00_3 <= D2_3;f01_3 <= d3_01;f02_3 <= d3_02;f03_3 <= d3_3;f10_3 <= d2_10;f20_3 <= d2_20;f30_3 <= d2_3;
                seq_4 <= ref[41:36];targ_4 <= read[53:48];f00_4 <= D3_3;f01_4 <= d4_01;f02_4 <= d4_02;f03_4 <= d4_3;f10_4 <= d3_10;f20_4 <= d3_20;f30_4 <= d3_3;     
                seq_5 <= ref[47:42];targ_5 <= read[47:42];f00_5 <= D4_3;f01_5 <= d5_01;f02_5 <= d5_02;f03_5 <= d5_3;f10_5 <= d4_10;f20_5 <= d4_20;f30_5 <= d4_3;
                seq_6 <= ref[53:48];targ_6 <= read[41:36];f00_6 <= D5_3;f01_6 <= d6_01;f02_6 <= d6_02;f03_6 <= d6_3;f10_6 <= d5_10;f20_6 <= d5_20;f30_6 <= d5_3;
                seq_7 <= ref[59:54];targ_7 <= read[35:30];f00_7 <= D6_3;f01_7 <= d7_01;f02_7 <= d7_02;f03_7 <= d7_3;f10_7 <= d6_10;f20_7 <= d6_20;f30_7 <= d6_3;
                seq_8 <= ref[65:60];targ_8 <= read[29:24];f00_8 <= D7_3;f01_8 <= d8_01;f02_8 <= d8_02;f03_8 <= d8_3;f10_8 <= d7_10;f20_8 <= d7_20;f30_8 <= d7_3;
                seq_9 <= ref[71:66];targ_9 <= read[23:18];f00_9 <= l;f01_9 <= l;f02_9 <= l;f03_9 <= l;f10_9 <= d8_10;f20_9 <= d8_20;f30_9 <= d8_3;
                state <= state + 1;
            end
       7'd28:
            begin
                seq_1 <= ref[17:12];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= d1_01;f02_1 <= d1_02;f03_1 <= d1_3;f10_1 <= l;f20_1 <= l;f30_1 <= l;
                seq_2 <= ref[23:18];targ_2 <= read[65:60];f00_2 <= D1_3;f01_2 <= d2_01;f02_2 <= d2_02;f03_2 <= d2_3;f10_2 <= d1_10;f20_2 <= d1_20;f30_2 <= d1_3;
                seq_3 <= ref[29:24];targ_3 <= read[59:54];f00_3 <= D2_3;f01_3 <= d3_01;f02_3 <= d3_02;f03_3 <= d3_3;f10_3 <= d2_10;f20_3 <= d2_20;f30_3 <= d2_3;
                seq_4 <= ref[35:30];targ_4 <= read[53:48];f00_4 <= D3_3;f01_4 <= d4_01;f02_4 <= d4_02;f03_4 <= d4_3;f10_4 <= d3_10;f20_4 <= d3_20;f30_4 <= d3_3;     
                seq_5 <= ref[41:36];targ_5 <= read[47:42];f00_5 <= D4_3;f01_5 <= d5_01;f02_5 <= d5_02;f03_5 <= d5_3;f10_5 <= d4_10;f20_5 <= d4_20;f30_5 <= d4_3;
                seq_6 <= ref[47:42];targ_6 <= read[41:36];f00_6 <= D5_3;f01_6 <= d6_01;f02_6 <= d6_02;f03_6 <= d6_3;f10_6 <= d5_10;f20_6 <= d5_20;f30_6 <= d5_3;
                seq_7 <= ref[53:48];targ_7 <= read[35:30];f00_7 <= D6_3;f01_7 <= d7_01;f02_7 <= d7_02;f03_7 <= d7_3;f10_7 <= d6_10;f20_7 <= d6_20;f30_7 <= d6_3;
                seq_8 <= ref[59:54];targ_8 <= read[29:24];f00_8 <= D7_3;f01_8 <= d8_01;f02_8 <= d8_02;f03_8 <= d8_3;f10_8 <= d7_10;f20_8 <= d7_20;f30_8 <= d7_3;
                seq_9 <= ref[65:60];targ_9 <= read[23:18];f00_9 <= D8_3;f01_9 <= d9_01;f02_9 <= d9_02;f03_9 <= d9_3;f10_9 <= d8_10;f20_9 <= d8_20;f30_9 <= d8_3;
                seq_10 <= ref[71:66];targ_10 <= read[17:12];f00_10 <= l;f01_10 <= l;f02_10 <= l;f03_10 <= l;f10_10 <= d9_10;f20_10 <= d9_20;f30_10 <= d9_3;
                state <= state + 1;
            end 
       7'd31:
            begin
                seq_1 <= ref[11:6];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= d1_01;f02_1 <= d1_02;f03_1 <= d1_3;f10_1 <= l;f20_1 <= l;f30_1 <= l;
                seq_2 <= ref[17:12];targ_2 <= read[65:60];f00_2 <= D1_3;f01_2 <= d2_01;f02_2 <= d2_02;f03_2 <= d2_3;f10_2 <= d1_10;f20_2 <= d1_20;f30_2 <= d1_3;
                seq_3 <= ref[23:18];targ_3 <= read[59:54];f00_3 <= D2_3;f01_3 <= d3_01;f02_3 <= d3_02;f03_3 <= d3_3;f10_3 <= d2_10;f20_3 <= d2_20;f30_3 <= d2_3;
                seq_4 <= ref[29:24];targ_4 <= read[53:48];f00_4 <= D3_3;f01_4 <= d4_01;f02_4 <= d4_02;f03_4 <= d4_3;f10_4 <= d3_10;f20_4 <= d3_20;f30_4 <= d3_3;     
                seq_5 <= ref[35:30];targ_5 <= read[47:42];f00_5 <= D4_3;f01_5 <= d5_01;f02_5 <= d5_02;f03_5 <= d5_3;f10_5 <= d4_10;f20_5 <= d4_20;f30_5 <= d4_3;
                seq_6 <= ref[41:36];targ_6 <= read[41:36];f00_6 <= D5_3;f01_6 <= d6_01;f02_6 <= d6_02;f03_6 <= d6_3;f10_6 <= d5_10;f20_6 <= d5_20;f30_6 <= d5_3;
                seq_7 <= ref[47:42];targ_7 <= read[35:30];f00_7 <= D6_3;f01_7 <= d7_01;f02_7 <= d7_02;f03_7 <= d7_3;f10_7 <= d6_10;f20_7 <= d6_20;f30_7 <= d6_3;
                seq_8 <= ref[53:48];targ_8 <= read[29:24];f00_8 <= D7_3;f01_8 <= d8_01;f02_8 <= d8_02;f03_8 <= d8_3;f10_8 <= d7_10;f20_8 <= d7_20;f30_8 <= d7_3;
                seq_9 <= ref[59:54];targ_9 <= read[23:18];f00_9 <= D8_3;f01_9 <= d9_01;f02_9 <= d9_02;f03_9 <= d9_3;f10_9 <= d8_10;f20_9 <= d8_20;f30_9 <= d8_3;
                seq_10 <= ref[65:60];targ_10 <= read[17:12];f00_10 <= D9_3;f01_10 <= d10_01;f02_10 <= d10_02;f03_10 <= d10_3;f10_10 <= d9_10;f20_10 <= d9_20;f30_10 <= d9_3;
                seq_11 <= ref[71:66];targ_11 <= read[11:6];f00_11 <= l;f01_11 <= l;f02_11 <= l;f03_11 <= l;f10_11 <= d10_10;f20_11 <= d10_20;f30_11 <= d10_3;
                state <= state + 1;
            end
       7'd34:
            begin
                seq_1 <= ref[5:0];targ_1 <= read[71:66];f00_1 <= l;f01_1 <= d1_01;f02_1 <= d1_02;f03_1 <= d1_3;f10_1 <= l;f20_1 <= l;f30_1 <= l;
                seq_2 <= ref[11:6];targ_2 <= read[65:60];f00_2 <= D1_3;f01_2 <= d2_01;f02_2 <= d2_02;f03_2 <= d2_3;f10_2 <= d1_10;f20_2 <= d1_20;f30_2 <= d1_3;
                seq_3 <= ref[17:12];targ_3 <= read[59:54];f00_3 <= D2_3;f01_3 <= d3_01;f02_3 <= d3_02;f03_3 <= d3_3;f10_3 <= d2_10;f20_3 <= d2_20;f30_3 <= d2_3;
                seq_4 <= ref[23:18];targ_4 <= read[53:48];f00_4 <= D3_3;f01_4 <= d4_01;f02_4 <= d4_02;f03_4 <= d4_3;f10_4 <= d3_10;f20_4 <= d3_20;f30_4 <= d3_3;     
                seq_5 <= ref[29:24];targ_5 <= read[47:42];f00_5 <= D4_3;f01_5 <= d5_01;f02_5 <= d5_02;f03_5 <= d5_3;f10_5 <= d4_10;f20_5 <= d4_20;f30_5 <= d4_3;
                seq_6 <= ref[35:30];targ_6 <= read[41:36];f00_6 <= D5_3;f01_6 <= d6_01;f02_6 <= d6_02;f03_6 <= d6_3;f10_6 <= d5_10;f20_6 <= d5_20;f30_6 <= d5_3;
                seq_7 <= ref[41:36];targ_7 <= read[35:30];f00_7 <= D6_3;f01_7 <= d7_01;f02_7 <= d7_02;f03_7 <= d7_3;f10_7 <= d6_10;f20_7 <= d6_20;f30_7 <= d6_3;
                seq_8 <= ref[47:42];targ_8 <= read[29:24];f00_8 <= D7_3;f01_8 <= d8_01;f02_8 <= d8_02;f03_8 <= d8_3;f10_8 <= d7_10;f20_8 <= d7_20;f30_8 <= d7_3;
                seq_9 <= ref[53:48];targ_9 <= read[23:18];f00_9 <= D8_3;f01_9 <= d9_01;f02_9 <= d9_02;f03_9 <= d9_3;f10_9 <= d8_10;f20_9 <= d8_20;f30_9 <= d8_3;
                seq_10 <= ref[59:54];targ_10 <= read[17:12];f00_10 <= D9_3;f01_10 <= d10_01;f02_10 <= d10_02;f03_10 <= d10_3;f10_10 <= d9_10;f20_10 <= d9_20;f30_10 <= d9_3;
                seq_11 <= ref[65:60];targ_11 <= read[11:6];f00_11 <= D10_3;f01_11 <= d11_01;f02_11 <= d11_02;f03_11 <= d11_3;f10_11 <= d10_10;f20_11 <= d10_20;f30_11 <= d10_3;
                seq_12 <= ref[71:66];targ_12 <= read[5:0];f00_12 <= l;f01_12 <= l;f02_12 <= l;f03_12 <= l;f10_12 <= d11_10;f20_12 <= d11_20;f30_12 <= d11_3;
                state <= state + 1;
            end    
      7'd37:
            begin
                seq_12 <= ref[5:0];targ_12 <= read[65:60];f00_12 <= D1_3;f01_12 <= d2_01;f02_12 <= d2_02;f03_12 <= d2_3;f10_12 <= d1_10;f20_12 <= d1_20;f30_12 <= d1_3;
                seq_11 <= ref[11:6];targ_11 <= read[59:54];f00_11 <= D2_3;f01_11 <= d3_01;f02_11 <= d3_02;f03_11 <= d3_3;f10_11 <= d2_10;f20_11 <= d2_20;f30_11 <= d2_3;
                seq_10 <= ref[17:12];targ_10 <= read[53:48];f00_10 <= D3_3;f01_10 <= d4_01;f02_10 <= d4_02;f03_10 <= d4_3;f10_10 <= d3_10;f20_10 <= d3_20;f30_10 <= d3_3;
                seq_9 <= ref[23:18];targ_9 <= read[47:42];f00_9 <= D4_3;f01_9 <= d5_01;f02_9 <= d5_02;f03_9 <= d5_3;f10_9 <= d4_10;f20_9 <= d4_20;f30_9 <= d4_3;     
                seq_8 <= ref[29:24];targ_8 <= read[41:36];f00_8 <= D5_3;f01_8 <= d6_01;f02_8 <= d6_02;f03_8 <= d6_3;f10_8 <= d5_10;f20_8 <= d5_20;f30_8 <= d5_3;
                seq_7 <= ref[35:30];targ_7 <= read[35:30];f00_7 <= D6_3;f01_7 <= d7_01;f02_7 <= d7_02;f03_7 <= d7_3;f10_7 <= d6_10;f20_7 <= d6_20;f30_7 <= d6_3;
                seq_6 <= ref[41:36];targ_6 <= read[29:24];f00_6 <= D7_3;f01_6 <= d8_01;f02_6 <= d8_02;f03_6 <= d8_3;f10_6 <= d7_10;f20_6 <= d7_20;f30_6 <= d7_3;
                seq_5 <= ref[47:42];targ_5 <= read[23:18];f00_5 <= D8_3;f01_5 <= d9_01;f02_5 <= d9_02;f03_5 <= d9_3;f10_5 <= d8_10;f20_5 <= d8_20;f30_5 <= d8_3;
                seq_4 <= ref[53:48];targ_4 <= read[17:12];f00_4 <= D9_3;f01_4 <= d10_01;f02_4 <= d10_02;f03_4 <= d10_3;f10_4 <= d9_10;f20_4 <= d9_20;f30_4 <= d9_3;
                seq_3 <= ref[59:54];targ_3 <= read[11:6];f00_3 <= D10_3;f01_3 <= d11_01;f02_3 <= d11_02;f03_3 <= d11_3;f10_3 <= d10_10;f20_3 <= d10_20;f30_3 <= d10_3;
                seq_2 <= ref[65:60];targ_2 <= read[5:0];f00_2 <= D11_3;f01_2 <= d12_01;f02_2 <= d12_02;f03_2 <= d12_3;f10_2 <= d11_10;f20_2 <= d11_20;f30_2 <= d11_3;
                state <= state + 1;
            end
     7'd40:
            begin
                seq_12 <= ref[5:0];targ_12 <= read[59:54];f00_12 <= D2_3;f01_12 <= d11_01;f02_12 <= d11_02;f03_12 <= d11_3;f10_12 <= d12_10;f20_12 <= d12_20;f30_12 <= d12_3;
                seq_11 <= ref[11:6];targ_11 <= read[53:48];f00_11 <= D3_3;f01_11 <= d10_01;f02_11 <= d10_02;f03_11 <= d10_3;f10_11 <= d11_10;f20_11 <= d11_20;f30_11 <= d11_3;
                seq_10 <= ref[17:12];targ_10 <= read[47:42];f00_10 <= D4_3;f01_10 <= d9_01;f02_10 <= d9_02;f03_10 <= d9_3;f10_10 <= d10_10;f20_10 <= d10_20;f30_10 <= d10_3;
                seq_9 <= ref[23:18];targ_9 <= read[41:36];f00_9 <= D5_3;f01_9 <= d8_01;f02_9 <= d8_02;f03_9 <= d8_3;f10_9 <= d9_10;f20_9 <= d9_20;f30_9 <= d9_3;     
                seq_8 <= ref[29:24];targ_8 <= read[35:30];f00_8 <= D6_3;f01_8 <= d7_01;f02_8 <= d7_02;f03_8 <= d7_3;f10_8 <= d8_10;f20_8 <= d8_20;f30_8 <= d8_3;
                seq_7 <= ref[35:30];targ_7 <= read[29:24];f00_7 <= D7_3;f01_7 <= d6_01;f02_7 <= d6_02;f03_7 <= d6_3;f10_7 <= d7_10;f20_7 <= d7_20;f30_7 <= d7_3;
                seq_6 <= ref[41:36];targ_6 <= read[23:18];f00_6 <= D8_3;f01_6 <= d5_01;f02_6 <= d5_02;f03_6 <= d5_3;f10_6 <= d6_10;f20_6 <= d6_20;f30_6 <= d6_3;
                seq_5 <= ref[47:42];targ_5 <= read[17:12];f00_5 <= D9_3;f01_5 <= d4_01;f02_5 <= d4_02;f03_5 <= d4_3;f10_5 <= d5_10;f20_5 <= d5_20;f30_5 <= d5_3;
                seq_4 <= ref[53:48];targ_4 <= read[11:6];f00_4 <= D10_3;f01_4 <= d3_01;f02_4 <= d3_02;f03_4 <= d3_3;f10_4 <= d4_10;f20_4 <= d4_20;f30_4 <= d4_3;
                seq_3 <= ref[59:54];targ_3 <= read[5:0];f00_3 <= D11_3;f01_3 <= d2_01;f02_3 <= d2_02;f03_3 <= d2_3;f10_3 <= d3_10;f20_3 <= d3_20;f30_3 <= d3_3;
                state <= state + 1;
            end
       7'd43:
            begin
                seq_12 <= ref[5:0];targ_12 <= read[53:48];f00_12 <= D11_3;f01_12 <= d11_01;f02_12 <= d11_02;f03_12 <= d11_3;f10_12 <= d12_10;f20_12 <= d12_20;f30_12 <= d12_3;
                seq_11 <= ref[11:6];targ_11 <= read[47:42];f00_11 <= D10_3;f01_11 <= d10_01;f02_11 <= d10_02;f03_11 <= d10_3;f10_11 <= d11_10;f20_11 <= d11_20;f30_11 <= d11_3;
                seq_10 <= ref[17:12];targ_10 <= read[41:36];f00_10 <= D9_3;f01_10 <= d9_01;f02_10 <= d9_02;f03_10 <= d9_3;f10_10 <= d10_10;f20_10 <= d10_20;f30_10 <= d10_3;
                seq_9 <= ref[23:18];targ_9 <= read[35:30];f00_9 <= D8_3;f01_9 <= d8_01;f02_9 <= d8_02;f03_9 <= d8_3;f10_9 <= d9_10;f20_9 <= d9_20;f30_9 <= d9_3;     
                seq_8 <= ref[29:24];targ_8 <= read[29:24];f00_8 <= D7_3;f01_8 <= d7_01;f02_8 <= d7_02;f03_8 <= d7_3;f10_8 <= d8_10;f20_8 <= d8_20;f30_8 <= d8_3;
                seq_7 <= ref[35:30];targ_7 <= read[23:18];f00_7 <= D6_3;f01_7 <= d6_01;f02_7 <= d6_02;f03_7 <= d6_3;f10_7 <= d7_10;f20_7 <= d7_20;f30_7 <= d7_3;
                seq_6 <= ref[41:36];targ_6 <= read[17:12];f00_6 <= D5_3;f01_6 <= d5_01;f02_6 <= d5_02;f03_6 <= d5_3;f10_6 <= d6_10;f20_6 <= d6_20;f30_6 <= d6_3;
                seq_5 <= ref[47:42];targ_5 <= read[11:6];f00_5 <= D4_3;f01_5 <= d4_01;f02_5 <= d4_02;f03_5 <= d4_3;f10_5 <= d5_10;f20_5 <= d5_20;f30_5 <= d5_3;
                seq_4 <= ref[53:48];targ_4 <= read[5:0];f00_4 <= D3_3;f01_4 <= d3_01;f02_4 <= d3_02;f03_4 <= d3_3;f10_4 <= d4_10;f20_4 <= d4_20;f30_4 <= d4_3;
                state <= state + 1;
            end
       7'd46:
            begin
                seq_12 <= ref[5:0];targ_12 <= read[47:42];f00_12 <= D11_3;f01_12 <= d11_01;f02_12 <= d11_02;f03_12 <= d11_3;f10_12 <= d12_10;f20_12 <= d12_20;f30_12 <= d12_3;
                seq_11 <= ref[11:6];targ_11 <= read[41:36];f00_11 <= D10_3;f01_11 <= d10_01;f02_11 <= d10_02;f03_11 <= d10_3;f10_11 <= d11_10;f20_11 <= d11_20;f30_11 <= d11_3;
                seq_10 <= ref[17:12];targ_10 <= read[35:30];f00_10 <= D9_3;f01_10 <= d9_01;f02_10 <= d9_02;f03_10 <= d9_3;f10_10 <= d10_10;f20_10 <= d10_20;f30_10 <= d10_3;
                seq_9 <= ref[23:18];targ_9 <= read[29:24];f00_9 <= D8_3;f01_9 <= d8_01;f02_9 <= d8_02;f03_9 <= d8_3;f10_9 <= d9_10;f20_9 <= d9_20;f30_9 <= d9_3;     
                seq_8 <= ref[29:24];targ_8 <= read[23:18];f00_8 <= D7_3;f01_8 <= d7_01;f02_8 <= d7_02;f03_8 <= d7_3;f10_8 <= d8_10;f20_8 <= d8_20;f30_8 <= d8_3;
                seq_7 <= ref[35:30];targ_7 <= read[17:12];f00_7 <= D6_3;f01_7 <= d6_01;f02_7 <= d6_02;f03_7 <= d6_3;f10_7 <= d7_10;f20_7 <= d7_20;f30_7 <= d7_3;
                seq_6 <= ref[41:36];targ_6 <= read[11:6];f00_6 <= D5_3;f01_6 <= d5_01;f02_6 <= d5_02;f03_6 <= d5_3;f10_6 <= d6_10;f20_6 <= d6_20;f30_6 <= d6_3;
                seq_5 <= ref[47:42];targ_5 <= read[5:0];f00_5 <= D4_3;f01_5 <= d4_01;f02_5 <= d4_02;f03_5 <= d4_3;f10_5 <= d5_10;f20_5 <= d5_20;f30_5 <= d5_3;
                state <= state + 1;
            end
       7'd49:
            begin
                seq_12 <= ref[5:0];targ_12 <= read[41:36];f00_12 <= D11_3;f01_12 <= d11_01;f02_12 <= d11_02;f03_12 <= d11_3;f10_12 <= d12_10;f20_12 <= d12_20;f30_12 <= d12_3;
                seq_11 <= ref[11:6];targ_11 <= read[35:30];f00_11 <= D10_3;f01_11 <= d10_01;f02_11 <= d10_02;f03_11 <= d10_3;f10_11 <= d11_10;f20_11 <= d11_20;f30_11 <= d11_3;
                seq_10 <= ref[17:12];targ_10 <= read[29:24];f00_10 <= D9_3;f01_10 <= d9_01;f02_10 <= d9_02;f03_10 <= d9_3;f10_10 <= d10_10;f20_10 <= d10_20;f30_10 <= d10_3;
                seq_9 <= ref[23:18];targ_9 <= read[23:18];f00_9 <= D8_3;f01_9 <= d8_01;f02_9 <= d8_02;f03_9 <= d8_3;f10_9 <= d9_10;f20_9 <= d9_20;f30_9 <= d9_3;     
                seq_8 <= ref[29:24];targ_8 <= read[17:12];f00_8 <= D7_3;f01_8 <= d7_01;f02_8 <= d7_02;f03_8 <= d7_3;f10_8 <= d8_10;f20_8 <= d8_20;f30_8 <= d8_3;
                seq_7 <= ref[35:30];targ_7 <= read[11:6];f00_7 <= D6_3;f01_7 <= d6_01;f02_7 <= d6_02;f03_7 <= d6_3;f10_7 <= d7_10;f20_7 <= d7_20;f30_7 <= d7_3;
                seq_6 <= ref[41:36];targ_6 <= read[5:0];f00_6 <= D5_3;f01_6 <= d5_01;f02_6 <= d5_02;f03_6 <= d5_3;f10_6 <= d6_10;f20_6 <= d6_20;f30_6 <= d6_3;
                state <= state + 1;
            end
       7'd52:
            begin
                seq_12 <= ref[5:0];targ_12 <= read[35:30];f00_12 <= D11_3;f01_12 <= d11_01;f02_12 <= d11_02;f03_12 <= d11_3;f10_12 <= d12_10;f20_12 <= d12_20;f30_12 <= d12_3;
                seq_11 <= ref[11:6];targ_11 <= read[29:24];f00_11 <= D10_3;f01_11 <= d10_01;f02_11 <= d10_02;f03_11 <= d10_3;f10_11 <= d11_10;f20_11 <= d11_20;f30_11 <= d11_3;
                seq_10 <= ref[17:12];targ_10 <= read[23:18];f00_10 <= D9_3;f01_10 <= d9_01;f02_10 <= d9_02;f03_10 <= d9_3;f10_10 <= d10_10;f20_10 <= d10_20;f30_10 <= d10_3;
                seq_9 <= ref[23:18];targ_9 <= read[17:12];f00_9 <= D8_3;f01_9 <= d8_01;f02_9 <= d8_02;f03_9 <= d8_3;f10_9 <= d9_10;f20_9 <= d9_20;f30_9 <= d9_3;     
                seq_8 <= ref[29:24];targ_8 <= read[11:6];f00_8 <= D7_3;f01_8 <= d7_01;f02_8 <= d7_02;f03_8 <= d7_3;f10_8 <= d8_10;f20_8 <= d8_20;f30_8 <= d8_3;
                seq_7 <= ref[35:30];targ_7 <= read[5:0];f00_7 <= D6_3;f01_7 <= d6_01;f02_7 <= d6_02;f03_7 <= d6_3;f10_7 <= d7_10;f20_7 <= d7_20;f30_7 <= d7_3;
                state <= state + 1;
            end
       7'd55:
            begin
                seq_12 <= ref[5:0];targ_12 <= read[29:24];f00_12 <= D11_3;f01_12 <= d11_01;f02_12 <= d11_02;f03_12 <= d11_3;f10_12 <= d12_10;f20_12 <= d12_20;f30_12 <= d12_3;
                seq_11 <= ref[11:6];targ_11 <= read[23:18];f00_11 <= D10_3;f01_11 <= d10_01;f02_11 <= d10_02;f03_11 <= d10_3;f10_11 <= d11_10;f20_11 <= d11_20;f30_11 <= d11_3;
                seq_10 <= ref[17:12];targ_10 <= read[17:12];f00_10 <= D9_3;f01_10 <= d9_01;f02_10 <= d9_02;f03_10 <= d9_3;f10_10 <= d10_10;f20_10 <= d10_20;f30_10 <= d10_3;
                seq_9 <= ref[23:18];targ_9 <= read[11:6];f00_9 <= D8_3;f01_9 <= d8_01;f02_9 <= d8_02;f03_9 <= d8_3;f10_9 <= d9_10;f20_9 <= d9_20;f30_9 <= d9_3;     
                seq_8 <= ref[29:24];targ_8 <= read[5:0];f00_8 <= D7_3;f01_8 <= d7_01;f02_8 <= d7_02;f03_8 <= d7_3;f10_8 <= d8_10;f20_8 <= d8_20;f30_8 <= d8_3;
                state <= state + 1;
                
            end
       7'd58:
            begin
                seq_12 <= ref[5:0];targ_12 <= read[23:18];f00_12 <= D11_3;f01_12 <= d11_01;f02_12 <= d11_02;f03_12 <= d11_3;f10_12 <= d12_10;f20_12 <= d12_20;f30_12 <= d12_3;
                seq_11 <= ref[11:6];targ_11 <= read[17:12];f00_11 <= D10_3;f01_11 <= d10_01;f02_11 <= d10_02;f03_11 <= d10_3;f10_11 <= d11_10;f20_11 <= d11_20;f30_11 <= d11_3;
                seq_10 <= ref[17:12];targ_10 <= read[11:6];f00_10 <= D9_3;f01_10 <= d9_01;f02_10 <= d9_02;f03_10 <= d9_3;f10_10 <= d10_10;f20_10 <= d10_20;f30_10 <= d10_3;
                seq_9 <= ref[23:18];targ_9 <= read[5:0];f00_9 <= D8_3;f01_9 <= d8_01;f02_9 <= d8_02;f03_9 <= d8_3;f10_9 <= d9_10;f20_9 <= d9_20;f30_9 <= d9_3;     
                state <= state + 1;
                
                max <= d10_3; 
            end
       7'd61:
            begin
                seq_12 <= ref[5:0];targ_12 <= read[17:12];f00_12 <= D11_3;f01_12 <= d11_01;f02_12 <= d11_02;f03_12 <= d11_3;f10_12 <= d12_10;f20_12 <= d12_20;f30_12 <= d12_3;
             //   seq_11 <= ref[11:6];targ_11 <= read[11:6];f00_11 <= D10_3;f01_11 <= d10_01;f02_11 <= d10_02;f03_11 <= d10_3;f10_11 <= d11_10;f20_11 <= d11_20;f30_11 <= d11_3;
                seq_10 <= ref[17:12];targ_10 <= read[5:0];f00_10 <= D9_3;f01_10 <= d9_01;f02_10 <= d9_02;f03_10 <= d9_3;f10_10 <= d10_10;f20_10 <= d10_20;f30_10 <= d10_3;
                state <= state + 1;
                sig <= 2'b01;
                if(d10_01 >= max && d10_01 >= d10_02 && d10_01 >= d10_3 && d10_01 >= d11_10 && d10_01 >= d11_20 && d10_01 >= d11_3 ) 
                    begin
                        max <= d10_01;
                        loc1[7] <= 1'b1;
                    end
                 if(d10_02 >= max && d10_02 >= d10_01 && d10_02 >= d10_3 && d10_02 >= d11_10 && d10_02 >= d11_20 && d10_02 >= d11_3) 
                    begin
                        max <= d10_02;
                        loc1[8] <= 1'b1;
                    end
                 if(d10_3 >= max && d10_3 >= d10_02 && d10_3 >= d10_01 && d10_3 >= d11_10 && d10_3 >= d11_20 && d10_3 >= d11_3) 
                    begin
                        max <= d10_3;
                        loc1[9] <= 1'b1;
                    end
                 if(d11_10 >= max && d11_10 >= d10_02 && d11_10 >= d10_3 && d11_10 >= d10_01 && d11_10 >= d11_20 && d11_10 >= d11_3) 
                    begin
                        max <= d11_10;
                        loc1[5] <= 1'b1;
                    end
                 if(d11_20 >= max && d11_20 >= d10_02 && d11_20 >= d10_3 && d11_20 >= d10_01 && d11_20 >= d11_10 && d11_20 >= d11_3) 
                    begin
                        max <= d11_20;
                        loc1[4] <= 1'b1;
                    end
                 if(d11_3 >= max && d11_3 >= d10_02 && d11_3 >= d10_3 && d11_3 >= d10_01 && d11_3 >= d11_20 && d11_3 >= d11_10) 
                    begin
                        max <= d11_3;
                        loc1[3] <= 1'b1;
                    end
                if(max >= d11_3 && max >= d10_02 && max >= d10_3 && max >= d10_01 && max >= d11_20 && max >= d11_10)
                    begin
                        loc1[6] <= 1'b1;
                    end
            end
     7'd64:
            begin
              state <= state + 1;
                if(d10_01 >= max && d10_01 >= d10_02 && d10_01 >= d10_3 && d10_01 >= d12_10 && d10_01 >= d12_20 && d10_01 >= d12_3) 
                    begin
                       if(d10_01 == max) sig <= 2'b11;
                       else sig <= 2'b10;
                        max <= d10_01;
                        loc2[10] <= 1'b1;
                    end
                if(d10_02 >= max && d10_02 >= d10_01 && d10_02 >= d10_3 && d10_02 >= d12_10 && d10_02 >= d12_20 && d10_02 >= d12_3) 
                    begin
                        if(d10_02 == max) sig <= 2'b11;
                        else sig <= 2'b10;
                        max <= d10_02;
                        loc2[11] <= 1'b1;
                    end
                if(d10_3 >= max && d10_3 >= d10_02 && d10_3 >= d10_01 && d10_3 >= d12_10 && d10_3 >= d12_20 && d10_3 >= d12_3) 
                    begin
                        if(d10_3 == max) sig <= 2'b11;
                        else sig <= 2'b10;
                        max <= d10_3;                        
                        loc2[12] <= 1'b1;
                    end
                if(d12_10 >= max && d12_10 >= d10_02 && d12_10 >= d10_3 && d12_10 >= d10_01 && d12_10 >= d12_20 && d12_10 >= d12_3) 
                    begin
                        if(d12_10 == max) sig <= 2'b11;
                        else sig <= 2'b10;
                        max <= d12_10;                        
                        loc2[2] <= 1'b1;
                    end
                if(d12_20 >= max && d12_20 >= d10_02 && d12_20 >= d10_3 && d12_20 >= d10_01 && d12_20 >= d12_10 && d12_20 >= d12_3) 
                    begin
                        if(d12_20 == max) sig <= 2'b11;
                        else sig <= 2'b10;
                        max <= d12_20;                        
                        loc2[1] <= 1'b1;
                    end
                if(d12_3 >= max && d12_3 >= d10_02 && d12_3 >= d10_3 && d12_3 >= d10_01 && d12_3 >= d12_20 && d12_3 >= d12_10) 
                    begin
                        if(d12_3 == max) sig <= 2'b11;
                        else sig <= 2'b10;
                        max <= d12_3;                        
                        loc2[0] <= 1'b1;
                    end
            end
     7'd65: begin
             finish <= 1;
             max <= max;
             loc1 <= loc1;
             loc2 <= loc2;
             sig <= sig; 
             //rst1 <= 0;
//             seq_1 <= 6'b000000;targ_1 <= 6'b111111;f00_1 <= l;f01_1 <= l;f02_1 <= l;f03_1 <= l;f10_1 <= l;f20_1 <= l;f30_1 <= l;
//                 seq_2 <= 6'b000000;targ_2 <= 6'b111111;f00_2 <= l;f01_2 <= l;f02_2 <= l;f03_2 <= l;f10_2 <= l;f20_2 <= l;f30_2 <= l;
//                 seq_3 <= 6'b000000;targ_3 <= 6'b111111;f00_3 <= l;f01_3 <= l;f02_3 <= l;f03_3 <= l;f10_3 <= l;f20_3 <= l;f30_3 <= l;
//                 seq_4 <= 6'b000000;targ_4 <= 6'b111111;f00_4 <= l;f01_4 <= l;f02_4 <= l;f03_4 <= l;f10_4 <= l;f20_4 <= l;f30_4 <= l;
//                 seq_5 <= 6'b000000;targ_5 <= 6'b111111;f00_5 <= l;f01_5 <= l;f02_5 <= l;f03_5 <= l;f10_5 <= l;f20_5 <= l;f30_5 <= l;
//                 seq_6 <= 6'b000000;targ_6 <= 6'b111111;f00_6 <= l;f01_6 <= l;f02_6 <= l;f03_6 <= l;f10_6 <= l;f20_6 <= l;f30_6 <= l;
//                 seq_7 <= 6'b000000;targ_7 <= 6'b111111;f00_7 <= l;f01_7 <= l;f02_7 <= l;f03_7 <= l;f10_7 <= l;f20_7 <= l;f30_7 <= l;
//                 seq_8 <= 6'b000000;targ_8 <= 6'b111111;f00_8 <= l;f01_8 <= l;f02_8 <= l;f03_8 <= l;f10_8 <= l;f20_8 <= l;f30_8 <= l;
//                 seq_9 <= 6'b000000;targ_9 <= 6'b111111;f00_9 <= l;f01_9 <= l;f02_9 <= l;f03_9 <= l;f10_9 <= l;f20_9 <= l;f30_9 <= l;
//                 seq_10 <= 6'b000000;targ_10 <= 6'b111111;f00_10 <= l;f01_10 <= l;f02_10 <= l;f03_10 <= l;f10_10 <= l;f20_10 <= l;f30_10 <= l;
//                 seq_11 <= 6'b000000;targ_11 <= 6'b111111;f00_11 <= l;f01_11 <= l;f02_11 <= l;f03_11 <= l;f10_11 <= l;f20_11 <= l;f30_11 <= l;
//                 seq_12 <= 6'b000000;targ_12 <= 6'b111111;f00_12 <= l;f01_12 <= l;f02_12 <= l;f03_12 <= l;f10_12 <= l;f20_12 <= l;f30_12 <= l;
                         
//                 D1_3 <= 0;
//                 D2_3 <= 0;
//                 D3_3 <= 0;
//                 D4_3 <= 0;
//                 D5_3 <= 0;
//                 D6_3 <= 0;
//                 D7_3 <= 0;
//                 D8_3 <= 0;
//                 D9_3 <= 0;
//                 D10_3 <= 0;
//                 D11_3 <= 0;
//                 D12_3 <= 0;
                 
//                 rst1 <= 0;
            end
     
      default:begin
            //finish <= 0;
            //rst1 <= 1;
            state <= state + 1;
            end 
       endcase             
    end
end

endmodule